module testbench ();



endmodule
